`define clock_gen(i) logic clock; initial begin forever begin clock = 0; #``i``; clock = 1; #``i``; end end