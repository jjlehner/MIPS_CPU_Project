module S_PC_Branch_Adder(	
	input	logic [31:0]	SRC_A , SRC_B,	
    input   logic [2:0]    ALUControl,
	output	logic [31:0]	ALU_Result
);
