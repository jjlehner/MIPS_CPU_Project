/* moduledoc



*/

module instruction_cache (
    input [31:0][31:0] raw_data
  );
  

endmodule