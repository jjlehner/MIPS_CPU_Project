module S_AND_2(
    input logic A,
    input logic B ,
    output logic Y
);

assign Y = A & B

endmodule