/* moduledoc



*/


module memory_controller (

  );

endmodule