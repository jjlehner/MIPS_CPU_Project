module Harvard_RAM(
	Harvard_Interface_RAM_side hv
);
endmodule

