module Adder
(
	input 	logic [31:0] a,b,
	output 	logic [31:0] z
);

assign z = a + b;

endmodule