module datapath (
    input clock, reset
  );



endmodule