/* moduledoc

*/

module address_decoder (
    input [31:0] read_address,
    input [31:0] write_address
  );
  

endmodule